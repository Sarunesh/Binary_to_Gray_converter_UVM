`include "uvm_pkg.sv"
import uvm_pkg::*;
`include "b2g_common.sv"
`include "b2g_intf.sv"
`include "b2g_tx.sv"
`include "b2g_seq_lib.sv"
`include "b2g_sequencer.sv"
`include "b2g_driver.sv"
`include "b2g_monitor.sv"
`include "b2g_subscriber.sv"
`include "b2g_agent.sv"
`include "b2g_sbd.sv"
`include "b2g_env.sv"
`include "test_lib.sv"
`include "bin_2_gray.v"
`include "top.sv"
