interface b2g_intf(input logic rst);
	logic [CODE_LENGTH-1:0] binary;
	logic [CODE_LENGTH-1:0] gray;
endinterface
