typedef uvm_sequencer#(b2g_tx) b2g_sequencer;
